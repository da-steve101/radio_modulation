`timescale 1ns / 1ps

module conv_lyr1_test
#(
) ();

   reg clk;
   reg rst;
   reg vld_in;
   reg [1:0][7:0] data_in [1:0];
   wire 	  vld_out;
   wire [127:0]   data_out [0:0];
   reg [8:0] 	  out_cntr;

   /*
    python code:
def ary_to_hex( x ):
  hex_str = ""
  for i in range( int( len(x) / 4 ) ):
    total = 0
    for j in range( 4 ):
      total += x[4*i + j] << ( 3 - j )
    hex_str += hex( total )[-1]
  return hex_str

# input_arys = [ np.array( [ i + 4, 0, i + 3, 0, i + 2, 0 ] ) for i in range( 32 ) ]
input_arys = [ np.array( [ 0, i + 2, 0, i + 3, 0, i + 4 ] ) for i in range( 32 ) ]
input_arys[0][1] = 0
res = [ list( reversed( 1*(np.matmul( w, lyr1_w ) >= lyr1_c) ) )  for w in input_arys ]
mp_res = [ [ a | b for a, b in zip( res[2*j], res[2*j+1] ) ] for j in range(16) ]
mp_hex = [ "256'h" + ary_to_hex( x ) for x in mp_res ]
", ".join( mp_hex )
   */
   wire [127:0]  expected_out [512] = { 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282b01254, 128'h025c4090403811700b2101a282b01254, 128'h025c4090407811700b2101a282b01254, 128'h025c4090407811700b2181a282b01254, 128'h025c4090407811700ba181a282b01254, 128'h02544090407811700ba181a282b01254, 128'h02544090407811700ba181a282b81254, 128'h0214c090407811700ba181a282b81254, 128'h0014c090407811700ba181a282b81254, 128'h0014c890407811700ba181a282b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700fa181a202381254, 128'h0014c890407811701fa181a202381254, 128'h0014c890407811701fa181a202381244, 128'h0014c890407811701ea381a602381244, 128'h0014c890407811701ea381a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381204, 128'h0014c891407811501ea3858602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c890407811710be1818682b91c14, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282b01254, 128'h025c4090403811700b2101a282b01254, 128'h025c4090407811700b2101a282b01254, 128'h025c4090407811700b2181a282b01254, 128'h025c4090407811700ba181a282b01254, 128'h02544090407811700ba181a282b01254, 128'h02544090407811700ba181a282b81254, 128'h0214c090407811700ba181a282b81254, 128'h0014c090407811700ba181a282b81254, 128'h0014c890407811700ba181a282b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700fa181a202381254, 128'h0014c890407811701fa181a202381254, 128'h0014c890407811701fa181a202381244, 128'h0014c890407811701ea381a602381244, 128'h0014c890407811701ea381a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381204, 128'h0014c891407811501ea3858602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c890407811710be1818682b91c14, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282b01254, 128'h025c4090403811700b2101a282b01254, 128'h025c4090407811700b2101a282b01254, 128'h025c4090407811700b2181a282b01254, 128'h025c4090407811700ba181a282b01254, 128'h02544090407811700ba181a282b01254, 128'h02544090407811700ba181a282b81254, 128'h0214c090407811700ba181a282b81254, 128'h0014c090407811700ba181a282b81254, 128'h0014c890407811700ba181a282b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700fa181a202381254, 128'h0014c890407811701fa181a202381254, 128'h0014c890407811701fa181a202381244, 128'h0014c890407811701ea381a602381244, 128'h0014c890407811701ea381a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381204, 128'h0014c891407811501ea3858602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c890407811710be1818682b91c14, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282b01254, 128'h025c4090403811700b2101a282b01254, 128'h025c4090407811700b2101a282b01254, 128'h025c4090407811700b2181a282b01254, 128'h025c4090407811700ba181a282b01254, 128'h02544090407811700ba181a282b01254, 128'h02544090407811700ba181a282b81254, 128'h0214c090407811700ba181a282b81254, 128'h0014c090407811700ba181a282b81254, 128'h0014c890407811700ba181a282b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700fa181a202381254, 128'h0014c890407811701fa181a202381254, 128'h0014c890407811701fa181a202381244, 128'h0014c890407811701ea381a602381244, 128'h0014c890407811701ea381a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381204, 128'h0014c891407811501ea3858602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c890407811710be1818682b91c14, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282b01254, 128'h025c4090403811700b2101a282b01254, 128'h025c4090407811700b2101a282b01254, 128'h025c4090407811700b2181a282b01254, 128'h025c4090407811700ba181a282b01254, 128'h02544090407811700ba181a282b01254, 128'h02544090407811700ba181a282b81254, 128'h0214c090407811700ba181a282b81254, 128'h0014c090407811700ba181a282b81254, 128'h0014c890407811700ba181a282b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700fa181a202381254, 128'h0014c890407811701fa181a202381254, 128'h0014c890407811701fa181a202381244, 128'h0014c890407811701ea381a602381244, 128'h0014c890407811701ea381a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381204, 128'h0014c891407811501ea3858602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c890407811710be1818682b91c14, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282b01254, 128'h025c4090403811700b2101a282b01254, 128'h025c4090407811700b2101a282b01254, 128'h025c4090407811700b2181a282b01254, 128'h025c4090407811700ba181a282b01254, 128'h02544090407811700ba181a282b01254, 128'h02544090407811700ba181a282b81254, 128'h0214c090407811700ba181a282b81254, 128'h0014c090407811700ba181a282b81254, 128'h0014c890407811700ba181a282b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700fa181a202381254, 128'h0014c890407811701fa181a202381254, 128'h0014c890407811701fa181a202381244, 128'h0014c890407811701ea381a602381244, 128'h0014c890407811701ea381a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381204, 128'h0014c891407811501ea3858602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c890407811710be1818682b91c14, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282b01254, 128'h025c4090403811700b2101a282b01254, 128'h025c4090407811700b2101a282b01254, 128'h025c4090407811700b2181a282b01254, 128'h025c4090407811700ba181a282b01254, 128'h02544090407811700ba181a282b01254, 128'h02544090407811700ba181a282b81254, 128'h0214c090407811700ba181a282b81254, 128'h0014c090407811700ba181a282b81254, 128'h0014c890407811700ba181a282b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700fa181a202381254, 128'h0014c890407811701fa181a202381254, 128'h0014c890407811701fa181a202381244, 128'h0014c890407811701ea381a602381244, 128'h0014c890407811701ea381a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381204, 128'h0014c891407811501ea3858602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c890407811710be1818682b91c14, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282b01254, 128'h025c4090403811700b2101a282b01254, 128'h025c4090407811700b2101a282b01254, 128'h025c4090407811700b2181a282b01254, 128'h025c4090407811700ba181a282b01254, 128'h02544090407811700ba181a282b01254, 128'h02544090407811700ba181a282b81254, 128'h0214c090407811700ba181a282b81254, 128'h0014c090407811700ba181a282b81254, 128'h0014c890407811700ba181a282b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700fa181a202381254, 128'h0014c890407811701fa181a202381254, 128'h0014c890407811701fa181a202381244, 128'h0014c890407811701ea381a602381244, 128'h0014c890407811701ea381a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381204, 128'h0014c891407811501ea3858602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c890407811710be1818682b91c14, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282b01254, 128'h025c4090403811700b2101a282b01254, 128'h025c4090407811700b2101a282b01254, 128'h025c4090407811700b2181a282b01254, 128'h025c4090407811700ba181a282b01254, 128'h02544090407811700ba181a282b01254, 128'h02544090407811700ba181a282b81254, 128'h0214c090407811700ba181a282b81254, 128'h0014c090407811700ba181a282b81254, 128'h0014c890407811700ba181a282b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700fa181a202381254, 128'h0014c890407811701fa181a202381254, 128'h0014c890407811701fa181a202381244, 128'h0014c890407811701ea381a602381244, 128'h0014c890407811701ea381a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381204, 128'h0014c891407811501ea3858602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c890407811710be1818682b91c14, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282b01254, 128'h025c4090403811700b2101a282b01254, 128'h025c4090407811700b2101a282b01254, 128'h025c4090407811700b2181a282b01254, 128'h025c4090407811700ba181a282b01254, 128'h02544090407811700ba181a282b01254, 128'h02544090407811700ba181a282b81254, 128'h0214c090407811700ba181a282b81254, 128'h0014c090407811700ba181a282b81254, 128'h0014c890407811700ba181a282b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700fa181a202381254, 128'h0014c890407811701fa181a202381254, 128'h0014c890407811701fa181a202381244, 128'h0014c890407811701ea381a602381244, 128'h0014c890407811701ea381a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381204, 128'h0014c891407811501ea3858602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c890407811710be1818682b91c14, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282b01254, 128'h025c4090403811700b2101a282b01254, 128'h025c4090407811700b2101a282b01254, 128'h025c4090407811700b2181a282b01254, 128'h025c4090407811700ba181a282b01254, 128'h02544090407811700ba181a282b01254, 128'h02544090407811700ba181a282b81254, 128'h0214c090407811700ba181a282b81254, 128'h0014c090407811700ba181a282b81254, 128'h0014c890407811700ba181a282b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700fa181a202381254, 128'h0014c890407811701fa181a202381254, 128'h0014c890407811701fa181a202381244, 128'h0014c890407811701ea381a602381244, 128'h0014c890407811701ea381a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381204, 128'h0014c891407811501ea3858602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c890407811710be1818682b91c14, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282b01254, 128'h025c4090403811700b2101a282b01254, 128'h025c4090407811700b2101a282b01254, 128'h025c4090407811700b2181a282b01254, 128'h025c4090407811700ba181a282b01254, 128'h02544090407811700ba181a282b01254, 128'h02544090407811700ba181a282b81254, 128'h0214c090407811700ba181a282b81254, 128'h0014c090407811700ba181a282b81254, 128'h0014c890407811700ba181a282b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700fa181a202381254, 128'h0014c890407811701fa181a202381254, 128'h0014c890407811701fa181a202381244, 128'h0014c890407811701ea381a602381244, 128'h0014c890407811701ea381a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381204, 128'h0014c891407811501ea3858602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c890407811710be1818682b91c14, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282b01254, 128'h025c4090403811700b2101a282b01254, 128'h025c4090407811700b2101a282b01254, 128'h025c4090407811700b2181a282b01254, 128'h025c4090407811700ba181a282b01254, 128'h02544090407811700ba181a282b01254, 128'h02544090407811700ba181a282b81254, 128'h0214c090407811700ba181a282b81254, 128'h0014c090407811700ba181a282b81254, 128'h0014c890407811700ba181a282b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700fa181a202381254, 128'h0014c890407811701fa181a202381254, 128'h0014c890407811701fa181a202381244, 128'h0014c890407811701ea381a602381244, 128'h0014c890407811701ea381a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381204, 128'h0014c891407811501ea3858602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c890407811710be1818682b91c14, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282b01254, 128'h025c4090403811700b2101a282b01254, 128'h025c4090407811700b2101a282b01254, 128'h025c4090407811700b2181a282b01254, 128'h025c4090407811700ba181a282b01254, 128'h02544090407811700ba181a282b01254, 128'h02544090407811700ba181a282b81254, 128'h0214c090407811700ba181a282b81254, 128'h0014c090407811700ba181a282b81254, 128'h0014c890407811700ba181a282b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700fa181a202381254, 128'h0014c890407811701fa181a202381254, 128'h0014c890407811701fa181a202381244, 128'h0014c890407811701ea381a602381244, 128'h0014c890407811701ea381a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381204, 128'h0014c891407811501ea3858602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c890407811710be1818682b91c14, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282b01254, 128'h025c4090403811700b2101a282b01254, 128'h025c4090407811700b2101a282b01254, 128'h025c4090407811700b2181a282b01254, 128'h025c4090407811700ba181a282b01254, 128'h02544090407811700ba181a282b01254, 128'h02544090407811700ba181a282b81254, 128'h0214c090407811700ba181a282b81254, 128'h0014c090407811700ba181a282b81254, 128'h0014c890407811700ba181a282b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700fa181a202381254, 128'h0014c890407811701fa181a202381254, 128'h0014c890407811701fa181a202381244, 128'h0014c890407811701ea381a602381244, 128'h0014c890407811701ea381a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381204, 128'h0014c891407811501ea3858602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c890407811710be1818682b91c14, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282b01254, 128'h025c4090403811700b2101a282b01254, 128'h025c4090407811700b2101a282b01254, 128'h025c4090407811700b2181a282b01254, 128'h025c4090407811700ba181a282b01254, 128'h02544090407811700ba181a282b01254, 128'h02544090407811700ba181a282b81254, 128'h0214c090407811700ba181a282b81254, 128'h0014c090407811700ba181a282b81254, 128'h0014c890407811700ba181a282b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700fa181a202381254, 128'h0014c890407811701fa181a202381254, 128'h0014c890407811701fa181a202381244, 128'h0014c890407811701ea381a602381244, 128'h0014c890407811701ea381a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381204, 128'h0014c891407811501ea3858602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c890407011710be1818682b91c14 };

always @( posedge clk ) begin
   if ( rst ) begin
      data_in[0] <= 16'h2;
      data_in[1] <= 16'h1;
      vld_in <= 0;
      out_cntr <= 0;
   end else begin
      vld_in <= 1;
      if ( vld_in ) begin
	 data_in[0] <= ( data_in[0] + 2 ) % 64;
	 data_in[1] <= ( data_in[1] + 2 ) % 64;
      end
      if ( vld_out ) begin
	 out_cntr <= out_cntr + 1;
	 if ( data_out[0] != expected_out[out_cntr % 512] ) begin
	    $display( "ASSERTION FAILED: data_out = %h, expected_out = %h", data_out[0], expected_out[out_cntr % 512] );
	 end
	 if ( out_cntr == 1500 ) begin
	    $finish;
	 end
      end
   end
end

lyr1 lyr1_inst
(
.clk(clk),
.rst(rst),
.vld_in(vld_in),
.data_in(data_in),
.vld_out(vld_out),
.data_out(data_out)
);

initial begin
   clk = 1;
   rst = 1;
   #10;
   rst = 0;
end

always begin
   #1;
   clk = !clk;
end

endmodule
