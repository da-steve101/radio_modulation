`timescale 1ns / 1ps

module conv_lyr2_test
#(
) ();

   reg clk;
   reg rst;
   reg vld_in;
   reg [255:0] data_in;
   wire 	  vld_out;
   wire [255:0]   data_out;
   reg [3:0] 	  out_cntr;
   reg [3:0] 	  in_cntr;

   /*
    python code:
def get_lyr( fname ):
  f = open( fname )
  rdr = csv.reader( f )
  return np.array( [ [ float(x) for x in y ] for y in rdr ] )

def ary_to_hex( x ):
  hex_str = ""
  for i in range( int( len(x) / 4 ) ):
    total = 0
    for j in range( 4 ):
      total += x[4*i + j] << ( 3 - j )
    hex_str += hex( total )[-1]
  return hex_str

def hex_to_ary( x ):
  all_bin = []
  for c in x:
    for b in format( int( c, 16 ), '004b' ):
      all_bin += [ int(b) ]
  return np.array( all_bin )

def hex_or( a, b ):
  hex_str = ""
  for x, y in zip( a, b ):
    hex_str += hex( int( x, 16 ) | int( y, 16 ) )[-1]
  return hex_str

def hex_xor( a, b ):
  hex_str = ""
  for x, y in zip( a, b ):
   hex_str += hex( int( x, 16 ) ^ int( y, 16 ) )[-1]
  return hex_str

lyr1_w = get_lyr( "vgg_conv_lyr_1.csv" )
lyr2_w = get_lyr( "vgg_conv_lyr_2.csv" )
f = open( "vgg_c_vec_lyr_1.csv" )
rdr = csv.reader( f )
lyr1_c = np.array( [ [ float(x) for x in y ] for y in rdr ] )
f = open( "vgg_c_vec_lyr_2.csv" )
rdr = csv.reader( f )
lyr2_c = np.array( [ [ float(x) for x in y ] for y in rdr ] )
lyr1_w = np.round( lyr1_w * ( 1 << 6 ) )
lyr1_c = lyr1_c * ( 1 << 6 )
input_arys = [ np.array( [ i + 4, 0, i + 3, 0, i + 2, 0 ] ) for i in range( 32 ) ]
input_arys[0][-2] = 0
res_1 = [ list( reversed( 1*(np.matmul( w, lyr1_w ) >= lyr1_c) ) )  for w in input_arys ]
mp_res = [ [ a | b for a, b in zip( res_1[2*j], res_1[2*j+1] ) ] for j in range(16) ]
input_arys = [ np.array( [ mp_res[i+1], mp_res[i], mp_res[i-1] ] ) for i in range( 15 ) ]
input_arys[0][-1] = 0*input_arys[0][-1]
input_arys = [ np.reshape( x, 3*256 ) for x in input_arys ]
res_2 = [ list( reversed( 1*(np.matmul( w, lyr2_w ) >= lyr2_c) ) )  for w in input_arys ]
mp_res = [ [ a | b for a, b in zip( res_2[2*j][0], res_2[2*j+1][0] ) ] for j in range(7) ]
mp_hex = [ "256'h" + ary_to_hex( x ) for x in mp_res ]
", ".join( mp_hex )
   */
   /*
   wire [255:0]   expected_in [16] = { 256'h0, 256'h0, 256'h0, 256'h0, 256'h0, 256'h0, 256'h0, 256'h0, 256'h0, 256'h0, 256'h0, 256'h0, 256'h0, 256'h0, 256'h0, 256'h0 };
   wire [255:0]   expected_out [7] = { 256'h89456bb09537410d56c038e2a8828061781420c8829c0b0d218088446a5dcd05, 256'h89456bb09537410d56c038e2a8828061781420c8829c0b0d218088446a5dcd05, 256'h89456bb09537410d56c038e2a8828061781420c8829c0b0d218088446a5dcd05, 256'h89456bb09537410d56c038e2a8828061781420c8829c0b0d218088446a5dcd05, 256'h89456bb09537410d56c038e2a8828061781420c8829c0b0d218088446a5dcd05, 256'h89456bb09537410d56c038e2a8828061781420c8829c0b0d218088446a5dcd05, 256'h89456bb09537410d56c038e2a8828061781420c8829c0b0d218088446a5dcd05 };
   // a0b3ba5622110184b0d039411304281e86014115471c036ab082eca90dd6a291
    */
   /*
   wire [255:0]   expected_in [16] = { 256'h0000000000000000000000000000000000000000000000000000000000000001, 256'h0000000000000000000000000000000000000000000000000000000000000002, 256'h0000000000000000000000000000000000000000000000000000000000000004, 256'h0000000000000000000000000000000000000000000000000000000000000008, 256'h0000000000000000000000000000000000000000000000000000000000000010, 256'h0000000000000000000000000000000000000000000000000000000000000020, 256'h0000000000000000000000000000000000000000000000000000000000000040, 256'h0000000000000000000000000000000000000000000000000000000000000080, 256'h0000000000000000000000000000000000000000000000000000000000000100, 256'h0000000000000000000000000000000000000000000000000000000000000200, 256'h0000000000000000000000000000000000000000000000000000000000000400, 256'h0000000000000000000000000000000000000000000000000000000000000800, 256'h0000000000000000000000000000000000000000000000000000000000001000, 256'h0000000000000000000000000000000000000000000000000000000000002000, 256'h0000000000000000000000000000000000000000000000000000000000004000, 256'h0000000000000000000000000000000000000000000000000000000000008000 };
   wire [255:0]   expected_out [7] = { 256'h89456bb09537410d56c338e2b8828061781420c8829c0b0d298088456a5dcd05, 256'h89456bb08537010d76c038e2a8828061781420ca829c0b0d218088456a5dcd45, 256'h89456bb09537410d56c238e2b8828061781420ca829c0b0d218088456a5dcd45, 256'h89456bb09537410d76c038e2a8828069781420ca809c0b0d298088446a5dcd55, 256'h89456bb09537410d76d038e2b8828061781420c8829c0b0d218088446a5dcd05, 256'h89456bb09537010d56c238e2a8828069781420ca829c0b0d298088446a5dcd05, 256'h89456bb09537410d56c238e2b8828061781420c8829c0b0d298088456a5dcd55 };
    */
   wire [255:0] expected_in [32] = { 256'h7640885406802bb16ca403d0a808310865a923002408db654888010108141699, 256'h7640885406802bb16c2403d0aa08310875a923002408d9654888010108541699, 256'h7640885406802bb16c2403d0aa08310c75a923002408d92548880101085c1699, 256'h7640885406802bb16c2403d0aa08310c75a923002408d92548880101085c1699, 256'h7640885406802bb16c240390aa08310c75a923002408d92548880101085c1699, 256'h7642885406002bb16c240390aa08310c75a923002408d92548880101085c1699, 256'h7642885416002bb16c240390aa08310c75a923002400d92548880101085c1699, 256'h7642885416002bb16c240390aa08310c75a923002400d92548880101085c1699, 256'h7642885416002bb16c240390aa08310c75a923002400d92548880101085c1699, 256'h7642885416002bb16c240390aa08310c75a923002400d92548880101085c1689, 256'h7642885416002bb02c240390aa08310c75a963002400d92548880101085c1689, 256'h7642885416002bb02c240390aa08310c75a963002400d92548880101085c1689, 256'h7642885416002bb02c240390aa08310c75a963002400d92548880101085c1689, 256'h7642885416002bb02c240390aa08310c75a973002400d92548880101085c1689, 256'h7642885516002bb02c240390aa08310475a973002400c92548880101085c1689, 256'h7642881516002bb03c240390aa28310455a973002400c92548888101085c1689, 256'h7642881516082bb034240390aa28310455a973002400c92548888101085c1689, 256'h7642881516082bb0342403908a28310455a973002400c92548888101085c1689, 256'h7642881516082bb0342403908a28310455a973002480c92548888101085c1689, 256'h7642881516082bb0342403908a28310455a973002480c92548898101085c1689, 256'h7642881516082bb0342403908a28310455a973002480c92548898101085c1689, 256'h7642881516082bb0342403908a28310454a973002480c92548898101085c16c9, 256'h7642880516082bb0342503908a28310454a973002480c92548898101085c16c9, 256'h7642880516082bb0342503908a28310454a973002480c92548898101085c16c9, 256'h7662080516082bb0346503908a28310454a973002480c92548898121085c16c9, 256'h7662080516082b30346502908a28310454a973002480c92548898121085c16c9, 256'h7662080516082330346512908a28310454a973002480c92548898121085c16c9, 256'h7662080516082330344512908a28310450a973002480c92548898121085c16c9, 256'h7662080516082330344512908a28310450a973002484c92548898121085c16c9, 256'h7662080516082330344512908a28310450a973002484c92508898121085c36c9, 256'h7663080516082370344512988a28310450a9f3002484c92528898121085c36c9, 256'h7663080516082370344512b88a20310450a9f3002484892528898121085c36c9 };

   wire [255:0] expected_out [16] = { 256'h7eb87bfce2ea30a27d60276dc8f8fdd2fedb5bbdbc22d0cf873da7c838876a13, 256'h7ef81a6ce2eb30a24d20274d49f8ddb2d6c9528dbc22d0cf973787ca3882aa30, 256'h7ef8184ce0eb34a24520254d49f855b2d7cb528ddc22d0cb973587c83882aa10, 256'h6ee8084ce0eb3422652025cd49f855b2d5cb528ddc22d0c31f7587c81082aa10, 256'h6ee80848e0eb3422652025cd49f855f2d5cbd28ddc22d2c31f7587c81082ea14, 256'h6e280a4ce2eb3420652025cd49f815f2d5cbd28dcc22c2d31b7587cc1082ea15, 256'hee280848e2eb34226520258d49f815f2d5cfd28dcca2c2d31b7187cc1082e815, 256'hee280848a5cb34226520258d49f015f2dd4fd28dc8a202d31971864c12c2e815, 256'hce280848e5c134206530208d48f015f29d47d28dc8a20283197386441282e805, 256'hce280848e5c134206530208d48f015f29d47d28cc8a20283197386441283e905, 256'hce2908c9e5c134206510208d49f015f29d47c28cc8a20283197386441283e905, 256'hce2908c9a5c135206710208d48d017e2bd47c28cc8aa0283997386441283e906, 256'h9c2948c9a5c135226790008f09d017e2bd47c2ac48aa0283996382443283ed07, 256'h982948c9a5c135267790288e09d017e2bf4783ac48aa0283196380453281cd06, 256'h982948c985c135266790288e09c007eabf4783ac48a8028119c3804532c1ed04, 256'h990149d9a5c137067710080e08c0046abb0783ac40a802a119c380450249cc04 };

always @( posedge clk ) begin
   if ( rst ) begin
      vld_in <= 0;
      out_cntr <= 0;
      in_cntr <= 0;
   end else begin
      vld_in <= 1;
      in_cntr <= in_cntr + 1;
      data_in <= expected_in[in_cntr];
      if ( vld_out ) begin
	 out_cntr <= out_cntr + 1;
	 if ( data_out != expected_out[out_cntr] ) begin
	    $display( "ASSERTION FAILED:\ndata_out     = %h\nexpected_out[%h] = %h", data_out, out_cntr, expected_out[out_cntr] );
	 end
	 if ( out_cntr == 6 ) begin
	    $finish;
	 end
      end
   end
end

lyr2 lyr2_inst
(
.clk(clk),
.rst(rst),
.vld_in(vld_in),
.data_in(data_in),
.vld_out(vld_out),
.data_out(data_out)
);

initial begin
   clk = 1;
   rst = 1;
   #10;
   rst = 0;
   #2000;
   $finish;
end

always begin
   #1;
   clk = !clk;
end

endmodule

