`timescale 1ns / 1ps

module conv_lyr2_test
#(
) ();

   reg clk;
   reg rst;
   reg vld_in;
   wire 	  vld_out;
   wire [127:0]   data_out;
   reg [7:0] 	  out_cntr;
   reg [8:0] 	  in_cntr;

   wire [127:0]  expected_in [512] = { 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282b01254, 128'h025c4090403811700b2101a282b01254, 128'h025c4090407811700b2101a282b01254, 128'h025c4090407811700b2181a282b01254, 128'h025c4090407811700ba181a282b01254, 128'h02544090407811700ba181a282b01254, 128'h02544090407811700ba181a282b81254, 128'h0214c090407811700ba181a282b81254, 128'h0014c090407811700ba181a282b81254, 128'h0014c890407811700ba181a282b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700fa181a202381254, 128'h0014c890407811701fa181a202381254, 128'h0014c890407811701fa181a202381244, 128'h0014c890407811701ea381a602381244, 128'h0014c890407811701ea381a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381204, 128'h0014c891407811501ea3858602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c890407811710be1818682b91c14, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282b01254, 128'h025c4090403811700b2101a282b01254, 128'h025c4090407811700b2101a282b01254, 128'h025c4090407811700b2181a282b01254, 128'h025c4090407811700ba181a282b01254, 128'h02544090407811700ba181a282b01254, 128'h02544090407811700ba181a282b81254, 128'h0214c090407811700ba181a282b81254, 128'h0014c090407811700ba181a282b81254, 128'h0014c890407811700ba181a282b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700fa181a202381254, 128'h0014c890407811701fa181a202381254, 128'h0014c890407811701fa181a202381244, 128'h0014c890407811701ea381a602381244, 128'h0014c890407811701ea381a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381204, 128'h0014c891407811501ea3858602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c890407811710be1818682b91c14, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282b01254, 128'h025c4090403811700b2101a282b01254, 128'h025c4090407811700b2101a282b01254, 128'h025c4090407811700b2181a282b01254, 128'h025c4090407811700ba181a282b01254, 128'h02544090407811700ba181a282b01254, 128'h02544090407811700ba181a282b81254, 128'h0214c090407811700ba181a282b81254, 128'h0014c090407811700ba181a282b81254, 128'h0014c890407811700ba181a282b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700fa181a202381254, 128'h0014c890407811701fa181a202381254, 128'h0014c890407811701fa181a202381244, 128'h0014c890407811701ea381a602381244, 128'h0014c890407811701ea381a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381204, 128'h0014c891407811501ea3858602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c890407811710be1818682b91c14, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282b01254, 128'h025c4090403811700b2101a282b01254, 128'h025c4090407811700b2101a282b01254, 128'h025c4090407811700b2181a282b01254, 128'h025c4090407811700ba181a282b01254, 128'h02544090407811700ba181a282b01254, 128'h02544090407811700ba181a282b81254, 128'h0214c090407811700ba181a282b81254, 128'h0014c090407811700ba181a282b81254, 128'h0014c890407811700ba181a282b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700fa181a202381254, 128'h0014c890407811701fa181a202381254, 128'h0014c890407811701fa181a202381244, 128'h0014c890407811701ea381a602381244, 128'h0014c890407811701ea381a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381204, 128'h0014c891407811501ea3858602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c890407811710be1818682b91c14, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282b01254, 128'h025c4090403811700b2101a282b01254, 128'h025c4090407811700b2101a282b01254, 128'h025c4090407811700b2181a282b01254, 128'h025c4090407811700ba181a282b01254, 128'h02544090407811700ba181a282b01254, 128'h02544090407811700ba181a282b81254, 128'h0214c090407811700ba181a282b81254, 128'h0014c090407811700ba181a282b81254, 128'h0014c890407811700ba181a282b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700fa181a202381254, 128'h0014c890407811701fa181a202381254, 128'h0014c890407811701fa181a202381244, 128'h0014c890407811701ea381a602381244, 128'h0014c890407811701ea381a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381204, 128'h0014c891407811501ea3858602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c890407811710be1818682b91c14, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282b01254, 128'h025c4090403811700b2101a282b01254, 128'h025c4090407811700b2101a282b01254, 128'h025c4090407811700b2181a282b01254, 128'h025c4090407811700ba181a282b01254, 128'h02544090407811700ba181a282b01254, 128'h02544090407811700ba181a282b81254, 128'h0214c090407811700ba181a282b81254, 128'h0014c090407811700ba181a282b81254, 128'h0014c890407811700ba181a282b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700fa181a202381254, 128'h0014c890407811701fa181a202381254, 128'h0014c890407811701fa181a202381244, 128'h0014c890407811701ea381a602381244, 128'h0014c890407811701ea381a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381204, 128'h0014c891407811501ea3858602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c890407811710be1818682b91c14, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282b01254, 128'h025c4090403811700b2101a282b01254, 128'h025c4090407811700b2101a282b01254, 128'h025c4090407811700b2181a282b01254, 128'h025c4090407811700ba181a282b01254, 128'h02544090407811700ba181a282b01254, 128'h02544090407811700ba181a282b81254, 128'h0214c090407811700ba181a282b81254, 128'h0014c090407811700ba181a282b81254, 128'h0014c890407811700ba181a282b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700fa181a202381254, 128'h0014c890407811701fa181a202381254, 128'h0014c890407811701fa181a202381244, 128'h0014c890407811701ea381a602381244, 128'h0014c890407811701ea381a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381204, 128'h0014c891407811501ea3858602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c890407811710be1818682b91c14, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282b01254, 128'h025c4090403811700b2101a282b01254, 128'h025c4090407811700b2101a282b01254, 128'h025c4090407811700b2181a282b01254, 128'h025c4090407811700ba181a282b01254, 128'h02544090407811700ba181a282b01254, 128'h02544090407811700ba181a282b81254, 128'h0214c090407811700ba181a282b81254, 128'h0014c090407811700ba181a282b81254, 128'h0014c890407811700ba181a282b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700fa181a202381254, 128'h0014c890407811701fa181a202381254, 128'h0014c890407811701fa181a202381244, 128'h0014c890407811701ea381a602381244, 128'h0014c890407811701ea381a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381204, 128'h0014c891407811501ea3858602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c890407811710be1818682b91c14, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282b01254, 128'h025c4090403811700b2101a282b01254, 128'h025c4090407811700b2101a282b01254, 128'h025c4090407811700b2181a282b01254, 128'h025c4090407811700ba181a282b01254, 128'h02544090407811700ba181a282b01254, 128'h02544090407811700ba181a282b81254, 128'h0214c090407811700ba181a282b81254, 128'h0014c090407811700ba181a282b81254, 128'h0014c890407811700ba181a282b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700fa181a202381254, 128'h0014c890407811701fa181a202381254, 128'h0014c890407811701fa181a202381244, 128'h0014c890407811701ea381a602381244, 128'h0014c890407811701ea381a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381204, 128'h0014c891407811501ea3858602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c890407811710be1818682b91c14, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282b01254, 128'h025c4090403811700b2101a282b01254, 128'h025c4090407811700b2101a282b01254, 128'h025c4090407811700b2181a282b01254, 128'h025c4090407811700ba181a282b01254, 128'h02544090407811700ba181a282b01254, 128'h02544090407811700ba181a282b81254, 128'h0214c090407811700ba181a282b81254, 128'h0014c090407811700ba181a282b81254, 128'h0014c890407811700ba181a282b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700fa181a202381254, 128'h0014c890407811701fa181a202381254, 128'h0014c890407811701fa181a202381244, 128'h0014c890407811701ea381a602381244, 128'h0014c890407811701ea381a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381204, 128'h0014c891407811501ea3858602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c890407811710be1818682b91c14, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282b01254, 128'h025c4090403811700b2101a282b01254, 128'h025c4090407811700b2101a282b01254, 128'h025c4090407811700b2181a282b01254, 128'h025c4090407811700ba181a282b01254, 128'h02544090407811700ba181a282b01254, 128'h02544090407811700ba181a282b81254, 128'h0214c090407811700ba181a282b81254, 128'h0014c090407811700ba181a282b81254, 128'h0014c890407811700ba181a282b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700fa181a202381254, 128'h0014c890407811701fa181a202381254, 128'h0014c890407811701fa181a202381244, 128'h0014c890407811701ea381a602381244, 128'h0014c890407811701ea381a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381204, 128'h0014c891407811501ea3858602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c890407811710be1818682b91c14, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282b01254, 128'h025c4090403811700b2101a282b01254, 128'h025c4090407811700b2101a282b01254, 128'h025c4090407811700b2181a282b01254, 128'h025c4090407811700ba181a282b01254, 128'h02544090407811700ba181a282b01254, 128'h02544090407811700ba181a282b81254, 128'h0214c090407811700ba181a282b81254, 128'h0014c090407811700ba181a282b81254, 128'h0014c890407811700ba181a282b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700fa181a202381254, 128'h0014c890407811701fa181a202381254, 128'h0014c890407811701fa181a202381244, 128'h0014c890407811701ea381a602381244, 128'h0014c890407811701ea381a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381204, 128'h0014c891407811501ea3858602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c890407811710be1818682b91c14, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282b01254, 128'h025c4090403811700b2101a282b01254, 128'h025c4090407811700b2101a282b01254, 128'h025c4090407811700b2181a282b01254, 128'h025c4090407811700ba181a282b01254, 128'h02544090407811700ba181a282b01254, 128'h02544090407811700ba181a282b81254, 128'h0214c090407811700ba181a282b81254, 128'h0014c090407811700ba181a282b81254, 128'h0014c890407811700ba181a282b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700fa181a202381254, 128'h0014c890407811701fa181a202381254, 128'h0014c890407811701fa181a202381244, 128'h0014c890407811701ea381a602381244, 128'h0014c890407811701ea381a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381204, 128'h0014c891407811501ea3858602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c890407811710be1818682b91c14, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282b01254, 128'h025c4090403811700b2101a282b01254, 128'h025c4090407811700b2101a282b01254, 128'h025c4090407811700b2181a282b01254, 128'h025c4090407811700ba181a282b01254, 128'h02544090407811700ba181a282b01254, 128'h02544090407811700ba181a282b81254, 128'h0214c090407811700ba181a282b81254, 128'h0014c090407811700ba181a282b81254, 128'h0014c890407811700ba181a282b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700fa181a202381254, 128'h0014c890407811701fa181a202381254, 128'h0014c890407811701fa181a202381244, 128'h0014c890407811701ea381a602381244, 128'h0014c890407811701ea381a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381204, 128'h0014c891407811501ea3858602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c890407811710be1818682b91c14, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282b01254, 128'h025c4090403811700b2101a282b01254, 128'h025c4090407811700b2101a282b01254, 128'h025c4090407811700b2181a282b01254, 128'h025c4090407811700ba181a282b01254, 128'h02544090407811700ba181a282b01254, 128'h02544090407811700ba181a282b81254, 128'h0214c090407811700ba181a282b81254, 128'h0014c090407811700ba181a282b81254, 128'h0014c890407811700ba181a282b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700fa181a202381254, 128'h0014c890407811701fa181a202381254, 128'h0014c890407811701fa181a202381244, 128'h0014c890407811701ea381a602381244, 128'h0014c890407811701ea381a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381204, 128'h0014c891407811501ea3858602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c890407811710be1818682b91c14, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282901254, 128'h025c4090403811700b0101a282b01254, 128'h025c4090403811700b2101a282b01254, 128'h025c4090407811700b2101a282b01254, 128'h025c4090407811700b2181a282b01254, 128'h025c4090407811700ba181a282b01254, 128'h02544090407811700ba181a282b01254, 128'h02544090407811700ba181a282b81254, 128'h0214c090407811700ba181a282b81254, 128'h0014c090407811700ba181a282b81254, 128'h0014c890407811700ba181a282b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202b81254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700ba181a202381254, 128'h0014c890407811700fa181a202381254, 128'h0014c890407811701fa181a202381254, 128'h0014c890407811701fa181a202381244, 128'h0014c890407811701ea381a602381244, 128'h0014c890407811701ea381a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea385a602381244, 128'h0014c891407811701ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381244, 128'h0014c891407811501ea3858602381204, 128'h0014c891407811501ea3858602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c891407811501ea3c58602391004, 128'h0014c890407011710be1818682b91c14 };

   wire [127:0] expected_out [256] = { 128'h095ab9292a04b32bcc830750d339f1d7, 128'h0d58b9a92a04932bcc810750d321f1d7, 128'h0d58b9a92a029329cc830710d341f1d7, 128'h0d58b12922028729d5860714d340f1d7, 128'h0d583109a282470155860714d344f197, 128'h2d58b009a382470155860284834c7197, 128'h2d5820018082470155860284834c7197, 128'h2d5820018082470155820284834c7197, 128'h2d5820018182430055820a84a30c7195, 128'h6d5c20018182430055820a84a34ce1dd, 128'h6d5c28019182630055822a84a34c61dd, 128'h655c28019182630071832a04a34e41dc, 128'h255c28019182630071822a04a34e41d8, 128'h255c28019182630071a32a04a34e41d8, 128'h255e28019180630051a32804a34e01c8, 128'h655a2809b8527321e1a32f86934d2d87, 128'h0d58b929ab06d32bdc810790d32df5d7, 128'h0d58b9a92a04932bcc810750d321f1d7, 128'h0d58b9a92a029329cc830710d341f1d7, 128'h0d58b12922028729d5860714d340f1d7, 128'h0d583109a282470155860714d344f197, 128'h2d58b009a382470155860284834c7197, 128'h2d5820018082470155860284834c7197, 128'h2d5820018082470155820284834c7197, 128'h2d5820018182430055820a84a30c7195, 128'h6d5c20018182430055820a84a34ce1dd, 128'h6d5c28019182630055822a84a34c61dd, 128'h655c28019182630071832a04a34e41dc, 128'h255c28019182630071822a04a34e41d8, 128'h255c28019182630071a32a04a34e41d8, 128'h255e28019180630051a32804a34e01c8, 128'h655a2809b8527321e1a32f86934d2d87, 128'h0d58b929ab06d32bdc810790d32df5d7, 128'h0d58b9a92a04932bcc810750d321f1d7, 128'h0d58b9a92a029329cc830710d341f1d7, 128'h0d58b12922028729d5860714d340f1d7, 128'h0d583109a282470155860714d344f197, 128'h2d58b009a382470155860284834c7197, 128'h2d5820018082470155860284834c7197, 128'h2d5820018082470155820284834c7197, 128'h2d5820018182430055820a84a30c7195, 128'h6d5c20018182430055820a84a34ce1dd, 128'h6d5c28019182630055822a84a34c61dd, 128'h655c28019182630071832a04a34e41dc, 128'h255c28019182630071822a04a34e41d8, 128'h255c28019182630071a32a04a34e41d8, 128'h255e28019180630051a32804a34e01c8, 128'h655a2809b8527321e1a32f86934d2d87, 128'h0d58b929ab06d32bdc810790d32df5d7, 128'h0d58b9a92a04932bcc810750d321f1d7, 128'h0d58b9a92a029329cc830710d341f1d7, 128'h0d58b12922028729d5860714d340f1d7, 128'h0d583109a282470155860714d344f197, 128'h2d58b009a382470155860284834c7197, 128'h2d5820018082470155860284834c7197, 128'h2d5820018082470155820284834c7197, 128'h2d5820018182430055820a84a30c7195, 128'h6d5c20018182430055820a84a34ce1dd, 128'h6d5c28019182630055822a84a34c61dd, 128'h655c28019182630071832a04a34e41dc, 128'h255c28019182630071822a04a34e41d8, 128'h255c28019182630071a32a04a34e41d8, 128'h255e28019180630051a32804a34e01c8, 128'h655a2809b8527321e1a32f86934d2d87, 128'h0d58b929ab06d32bdc810790d32df5d7, 128'h0d58b9a92a04932bcc810750d321f1d7, 128'h0d58b9a92a029329cc830710d341f1d7, 128'h0d58b12922028729d5860714d340f1d7, 128'h0d583109a282470155860714d344f197, 128'h2d58b009a382470155860284834c7197, 128'h2d5820018082470155860284834c7197, 128'h2d5820018082470155820284834c7197, 128'h2d5820018182430055820a84a30c7195, 128'h6d5c20018182430055820a84a34ce1dd, 128'h6d5c28019182630055822a84a34c61dd, 128'h655c28019182630071832a04a34e41dc, 128'h255c28019182630071822a04a34e41d8, 128'h255c28019182630071a32a04a34e41d8, 128'h255e28019180630051a32804a34e01c8, 128'h655a2809b8527321e1a32f86934d2d87, 128'h0d58b929ab06d32bdc810790d32df5d7, 128'h0d58b9a92a04932bcc810750d321f1d7, 128'h0d58b9a92a029329cc830710d341f1d7, 128'h0d58b12922028729d5860714d340f1d7, 128'h0d583109a282470155860714d344f197, 128'h2d58b009a382470155860284834c7197, 128'h2d5820018082470155860284834c7197, 128'h2d5820018082470155820284834c7197, 128'h2d5820018182430055820a84a30c7195, 128'h6d5c20018182430055820a84a34ce1dd, 128'h6d5c28019182630055822a84a34c61dd, 128'h655c28019182630071832a04a34e41dc, 128'h255c28019182630071822a04a34e41d8, 128'h255c28019182630071a32a04a34e41d8, 128'h255e28019180630051a32804a34e01c8, 128'h655a2809b8527321e1a32f86934d2d87, 128'h0d58b929ab06d32bdc810790d32df5d7, 128'h0d58b9a92a04932bcc810750d321f1d7, 128'h0d58b9a92a029329cc830710d341f1d7, 128'h0d58b12922028729d5860714d340f1d7, 128'h0d583109a282470155860714d344f197, 128'h2d58b009a382470155860284834c7197, 128'h2d5820018082470155860284834c7197, 128'h2d5820018082470155820284834c7197, 128'h2d5820018182430055820a84a30c7195, 128'h6d5c20018182430055820a84a34ce1dd, 128'h6d5c28019182630055822a84a34c61dd, 128'h655c28019182630071832a04a34e41dc, 128'h255c28019182630071822a04a34e41d8, 128'h255c28019182630071a32a04a34e41d8, 128'h255e28019180630051a32804a34e01c8, 128'h655a2809b8527321e1a32f86934d2d87, 128'h0d58b929ab06d32bdc810790d32df5d7, 128'h0d58b9a92a04932bcc810750d321f1d7, 128'h0d58b9a92a029329cc830710d341f1d7, 128'h0d58b12922028729d5860714d340f1d7, 128'h0d583109a282470155860714d344f197, 128'h2d58b009a382470155860284834c7197, 128'h2d5820018082470155860284834c7197, 128'h2d5820018082470155820284834c7197, 128'h2d5820018182430055820a84a30c7195, 128'h6d5c20018182430055820a84a34ce1dd, 128'h6d5c28019182630055822a84a34c61dd, 128'h655c28019182630071832a04a34e41dc, 128'h255c28019182630071822a04a34e41d8, 128'h255c28019182630071a32a04a34e41d8, 128'h255e28019180630051a32804a34e01c8, 128'h655a2809b8527321e1a32f86934d2d87, 128'h0d58b929ab06d32bdc810790d32df5d7, 128'h0d58b9a92a04932bcc810750d321f1d7, 128'h0d58b9a92a029329cc830710d341f1d7, 128'h0d58b12922028729d5860714d340f1d7, 128'h0d583109a282470155860714d344f197, 128'h2d58b009a382470155860284834c7197, 128'h2d5820018082470155860284834c7197, 128'h2d5820018082470155820284834c7197, 128'h2d5820018182430055820a84a30c7195, 128'h6d5c20018182430055820a84a34ce1dd, 128'h6d5c28019182630055822a84a34c61dd, 128'h655c28019182630071832a04a34e41dc, 128'h255c28019182630071822a04a34e41d8, 128'h255c28019182630071a32a04a34e41d8, 128'h255e28019180630051a32804a34e01c8, 128'h655a2809b8527321e1a32f86934d2d87, 128'h0d58b929ab06d32bdc810790d32df5d7, 128'h0d58b9a92a04932bcc810750d321f1d7, 128'h0d58b9a92a029329cc830710d341f1d7, 128'h0d58b12922028729d5860714d340f1d7, 128'h0d583109a282470155860714d344f197, 128'h2d58b009a382470155860284834c7197, 128'h2d5820018082470155860284834c7197, 128'h2d5820018082470155820284834c7197, 128'h2d5820018182430055820a84a30c7195, 128'h6d5c20018182430055820a84a34ce1dd, 128'h6d5c28019182630055822a84a34c61dd, 128'h655c28019182630071832a04a34e41dc, 128'h255c28019182630071822a04a34e41d8, 128'h255c28019182630071a32a04a34e41d8, 128'h255e28019180630051a32804a34e01c8, 128'h655a2809b8527321e1a32f86934d2d87, 128'h0d58b929ab06d32bdc810790d32df5d7, 128'h0d58b9a92a04932bcc810750d321f1d7, 128'h0d58b9a92a029329cc830710d341f1d7, 128'h0d58b12922028729d5860714d340f1d7, 128'h0d583109a282470155860714d344f197, 128'h2d58b009a382470155860284834c7197, 128'h2d5820018082470155860284834c7197, 128'h2d5820018082470155820284834c7197, 128'h2d5820018182430055820a84a30c7195, 128'h6d5c20018182430055820a84a34ce1dd, 128'h6d5c28019182630055822a84a34c61dd, 128'h655c28019182630071832a04a34e41dc, 128'h255c28019182630071822a04a34e41d8, 128'h255c28019182630071a32a04a34e41d8, 128'h255e28019180630051a32804a34e01c8, 128'h655a2809b8527321e1a32f86934d2d87, 128'h0d58b929ab06d32bdc810790d32df5d7, 128'h0d58b9a92a04932bcc810750d321f1d7, 128'h0d58b9a92a029329cc830710d341f1d7, 128'h0d58b12922028729d5860714d340f1d7, 128'h0d583109a282470155860714d344f197, 128'h2d58b009a382470155860284834c7197, 128'h2d5820018082470155860284834c7197, 128'h2d5820018082470155820284834c7197, 128'h2d5820018182430055820a84a30c7195, 128'h6d5c20018182430055820a84a34ce1dd, 128'h6d5c28019182630055822a84a34c61dd, 128'h655c28019182630071832a04a34e41dc, 128'h255c28019182630071822a04a34e41d8, 128'h255c28019182630071a32a04a34e41d8, 128'h255e28019180630051a32804a34e01c8, 128'h655a2809b8527321e1a32f86934d2d87, 128'h0d58b929ab06d32bdc810790d32df5d7, 128'h0d58b9a92a04932bcc810750d321f1d7, 128'h0d58b9a92a029329cc830710d341f1d7, 128'h0d58b12922028729d5860714d340f1d7, 128'h0d583109a282470155860714d344f197, 128'h2d58b009a382470155860284834c7197, 128'h2d5820018082470155860284834c7197, 128'h2d5820018082470155820284834c7197, 128'h2d5820018182430055820a84a30c7195, 128'h6d5c20018182430055820a84a34ce1dd, 128'h6d5c28019182630055822a84a34c61dd, 128'h655c28019182630071832a04a34e41dc, 128'h255c28019182630071822a04a34e41d8, 128'h255c28019182630071a32a04a34e41d8, 128'h255e28019180630051a32804a34e01c8, 128'h655a2809b8527321e1a32f86934d2d87, 128'h0d58b929ab06d32bdc810790d32df5d7, 128'h0d58b9a92a04932bcc810750d321f1d7, 128'h0d58b9a92a029329cc830710d341f1d7, 128'h0d58b12922028729d5860714d340f1d7, 128'h0d583109a282470155860714d344f197, 128'h2d58b009a382470155860284834c7197, 128'h2d5820018082470155860284834c7197, 128'h2d5820018082470155820284834c7197, 128'h2d5820018182430055820a84a30c7195, 128'h6d5c20018182430055820a84a34ce1dd, 128'h6d5c28019182630055822a84a34c61dd, 128'h655c28019182630071832a04a34e41dc, 128'h255c28019182630071822a04a34e41d8, 128'h255c28019182630071a32a04a34e41d8, 128'h255e28019180630051a32804a34e01c8, 128'h655a2809b8527321e1a32f86934d2d87, 128'h0d58b929ab06d32bdc810790d32df5d7, 128'h0d58b9a92a04932bcc810750d321f1d7, 128'h0d58b9a92a029329cc830710d341f1d7, 128'h0d58b12922028729d5860714d340f1d7, 128'h0d583109a282470155860714d344f197, 128'h2d58b009a382470155860284834c7197, 128'h2d5820018082470155860284834c7197, 128'h2d5820018082470155820284834c7197, 128'h2d5820018182430055820a84a30c7195, 128'h6d5c20018182430055820a84a34ce1dd, 128'h6d5c28019182630055822a84a34c61dd, 128'h655c28019182630071832a04a34e41dc, 128'h255c28019182630071822a04a34e41d8, 128'h255c28019182630071a32a04a34e41d8, 128'h255e28019180630051a32804a34e01c8, 128'h655a2809b8527321e1a32f86934d2d87, 128'h0d58b929ab06d32bdc810790d32df5d7, 128'h0d58b9a92a04932bcc810750d321f1d7, 128'h0d58b9a92a029329cc830710d341f1d7, 128'h0d58b12922028729d5860714d340f1d7, 128'h0d583109a282470155860714d344f197, 128'h2d58b009a382470155860284834c7197, 128'h2d5820018082470155860284834c7197, 128'h2d5820018082470155820284834c7197, 128'h2d5820018182430055820a84a30c7195, 128'h6d5c20018182430055820a84a34ce1dd, 128'h6d5c28019182630055822a84a34c61dd, 128'h655c28019182630071832a04a34e41dc, 128'h255c28019182630071822a04a34e41d8, 128'h255c28019182630071a32a04a34e41d8, 128'h255e28019180630051a32804a34e01c8, 128'h6dde68499d52772029a32f86074d01e5 };

always @( posedge clk ) begin
   if ( rst ) begin
      vld_in <= 0;
      out_cntr <= 0;
      in_cntr <= 0;
   end else begin
      vld_in <= !vld_in;
      if ( vld_in ) begin
	 in_cntr <= in_cntr + 1;
      end
      if ( vld_out ) begin
	 out_cntr <= out_cntr + 1;
	 if ( data_out != expected_out[out_cntr % 256] ) begin
	    $display( "ASSERTION FAILED: data_out = %h, expected_out[%d] = %h", data_out, out_cntr, expected_out[out_cntr % 256] );
	 end
	 if ( out_cntr == 700 ) begin
	    $finish;
	 end
      end
   end
end

lyr2 lyr2_inst
(
.clk(clk),
.rst(rst),
.vld_in(vld_in),
.data_in(expected_in[in_cntr]),
.vld_out(vld_out),
.data_out(data_out)
);

initial begin
   clk = 1;
   rst = 1;
   #10;
   rst = 0;
   #2000;
   $finish;
end

always begin
   #1;
   clk = !clk;
end

endmodule

